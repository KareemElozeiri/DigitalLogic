module test_stopwatch();

logic clk,reset,enable,up;
logic[3:0] q0,q1,q2,q3;
stopwatch c(clk,up,enable,reset,q0,q1,q2,q3);
always #50 clk= ~clk;

initial begin
clk = 0;
reset = 1;
enable = 0;
up = 1;
#200;
reset = 1;
enable = 0;
up = 1;
#200;
reset = 1;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 0;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 1;
#200;
reset = 1;
enable = 1;
up = 1;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
reset = 0;
enable = 1;
up = 0;
#200;
$stop;
end 

endmodule 