module test_counter();
logic clk,reset,enable,up,load;
logic[3:0] load_signal;
logic[3:0] q;
logic next_counter_clk;
counter5 c(clk,reset,enable,up,load,load_signal,q,next_counter_clk);
always #50 clk= ~clk;

initial begin
clk = 0;
reset = 1;
enable = 0;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 1;
enable = 0;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 1;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 1;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 0;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 1;
enable = 1;
up = 1;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
reset = 0;
enable = 1;
up = 0;
load = 0;
load_signal = 4'b0011;
#200;
$stop;
end 

endmodule